float Mesh2_face_Stroemungsgeschwindigkeit_x_2d(nMesh2_data_time, nMesh2_layer_2d, nMesh2_face) ;
    Mesh2_face_Stroemungsgeschwindigkeit_x_2d:long_name = "Stroemungsgeschwindigkeit (x-Komponente), Face (Polygon)" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_x_2d:units = "m s-1" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_x_2d:name_id = 2 ; 
    Mesh2_face_Stroemungsgeschwindigkeit_x_2d:_FillValue = 1.e+31f ; 
    Mesh2_face_Stroemungsgeschwindigkeit_x_2d:cell_methods = "nMesh2_data_time: point nMesh2_layer_2d: mean area: point" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_x_2d:coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat Mesh2_face_z_face_2d" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_x_2d:grid_mapping = "Mesh2_crs" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_x_2d:standard_name = "sea_water_x_velocity" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_x_2d:mesh = "Mesh2" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_x_2d:location = "face" ; 
//    Mesh2_face_Stroemungsgeschwindigkeit_x_2d:davit_role = "visualization_variable" ;



float Mesh2_face_Stroemungsgeschwindigkeit_y_2d(nMesh2_data_time, nMesh2_layer_2d, nMesh2_face) ;
    Mesh2_face_Stroemungsgeschwindigkeit_y_2d:long_name = "Stroemungsgeschwindigkeit (y-Komponente), Face (Polygon)" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_y_2d:units = "m s-1" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_y_2d:name_id = 2 ; 
    Mesh2_face_Stroemungsgeschwindigkeit_y_2d:_FillValue = 1.e+31f ; 
    Mesh2_face_Stroemungsgeschwindigkeit_y_2d:cell_methods = "nMesh2_data_time: point nMesh2_layer_2d: mean area: point" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_y_2d:coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat Mesh2_face_z_face_2d" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_y_2d:grid_mapping = "Mesh2_crs" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_y_2d:standard_name = "sea_water_y_velocity" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_y_2d:mesh = "Mesh2" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_y_2d:location = "face" ; 
//    Mesh2_face_Stroemungsgeschwindigkeit_y_2d:davit_role = "visualization_variable" ;


float Mesh2_face_Stroemungsgeschwindigkeit_m_2d(nMesh2_data_time, nMesh2_layer_2d, nMesh2_face) ;
    Mesh2_face_Stroemungsgeschwindigkeit_m_2d:long_name = "Stroemungsgeschwindigkeit (Betrag), Face (Polygon)" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_m_2d:units = "m s-1" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_m_2d:name_id = 2 ; 
    Mesh2_face_Stroemungsgeschwindigkeit_m_2d:_FillValue = 1.e+31f ; 
    Mesh2_face_Stroemungsgeschwindigkeit_m_2d:cell_methods = "nMesh2_data_time: point nMesh2_layer_2d: mean area: point" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_m_2d:coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat Mesh2_face_z_face_2d" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_m_2d:grid_mapping = "Mesh2_crs" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_m_2d:standard_name = "magnitude_of_sea_water_velocity" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_m_2d:mesh = "Mesh2" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_m_2d:location = "face" ; 
//    Mesh2_face_Stroemungsgeschwindigkeit_m_2d:davit_role = "visualization_variable" ;

   
float Mesh2_face_Temperatur_3d(nMesh2_data_time, nMesh2_layer_3d, nMesh2_face) ;
    Mesh2_face_Temperatur_3d:long_name = "Temperatur, Face (Polygon)" ;
    Mesh2_face_Temperatur_3d:units = "degC" ;
    Mesh2_face_Temperatur_3d:name_id = 6 ;
    Mesh2_face_Temperatur_3d:_FillValue = 1.e+31f ;
    Mesh2_face_Temperatur_3d:cell_measures = "area: Mesh2_face_wet_area" ;
    Mesh2_face_Temperatur_3d:cell_methods = "nMesh2_data_time: point nMesh2_layer_3d: mean area: point" ;
    Mesh2_face_Temperatur_3d:coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat Mesh2_face_z_face_3d" ;
    Mesh2_face_Temperatur_3d:grid_mapping = "Mesh2_crs" ;
    Mesh2_face_Temperatur_3d:standard_name = "temperature" ;
    Mesh2_face_Temperatur_3d:mesh = "Mesh2" ;
    Mesh2_face_Temperatur_3d:location = "face" ;
//    Mesh2_face_Temperatur_3d:davit_role = "visualization_variable" ;

double Mesh2_face_depth_2d(nMesh2_time, nMesh2_face) ;
    Mesh2_face_depth_2d:long_name = "Topographie" ;
    Mesh2_face_depth_2d:units = "m" ;
    Mesh2_face_depth_2d:name_id = 17 ;
    Mesh2_face_depth_2d:valid_range = -8848., 11034. ;
    Mesh2_face_depth_2d:_FillValue = 1.e+31 ;
    Mesh2_face_depth_2d:cell_measures = "area: Mesh2_face_area" ;
    Mesh2_face_depth_2d:cell_methods = "nMesh2_time: mean area: mean" ;
    Mesh2_face_depth_2d:coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ;
    Mesh2_face_depth_2d:grid_mapping = "Mesh2_crs" ;
    Mesh2_face_depth_2d:standard_name = "sea_floor_depth_below_geoid" ;
    Mesh2_face_depth_2d:mesh = "Mesh2" ;
    Mesh2_face_depth_2d:location = "face" ;
//    Mesh2_face_depth_2d:davit_role = "visualization_variable" ;

float Mesh2_face_Wasserstand_2d(nMesh2_data_time, nMesh2_face) ;
    Mesh2_face_Wasserstand_2d:long_name = "Wasserstand, Face (Polygon)" ; 
    Mesh2_face_Wasserstand_2d:units = "m" ; 
    Mesh2_face_Wasserstand_2d:name_id = 3 ; 
    Mesh2_face_Wasserstand_2d:_FillValue = 1.e+31f ; 
    Mesh2_face_Wasserstand_2d:cell_measures = "area: Mesh2_face_wet_area" ; 
    Mesh2_face_Wasserstand_2d:cell_methods = "nMesh2_data_time: point area: mean" ; 
    Mesh2_face_Wasserstand_2d:coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ; 
    Mesh2_face_Wasserstand_2d:grid_mapping = "Mesh2_crs" ; 
    Mesh2_face_Wasserstand_2d:standard_name = "sea_surface_height" ; 
    Mesh2_face_Wasserstand_2d:mesh = "Mesh2" ; 
    Mesh2_face_Wasserstand_2d:location = "face" ; 

float Mesh2_face_Gesamtwassertiefe_2d(nMesh2_data_time, nMesh2_face) ;
    Mesh2_face_Gesamtwassertiefe_2d:long_name = "Gesamtwassertiefe [ face ]" ;
    Mesh2_face_Gesamtwassertiefe_2d:units = "m" ;
    Mesh2_face_Gesamtwassertiefe_2d:name_id = 16 ;
    Mesh2_face_Gesamtwassertiefe_2d:_FillValue = 1.e+31f ;
    Mesh2_face_Gesamtwassertiefe_2d:cell_methods = "nMesh2_data_time: point nMesh2_face: mean" ;
    Mesh2_face_Gesamtwassertiefe_2d:coordinates = "Mesh2_face_lon Mesh2_face_lat Mesh2_face_x Mesh2_face_y" ;
    Mesh2_face_Gesamtwassertiefe_2d:grid_mapping = "Mesh2_crs" ;
    Mesh2_face_Gesamtwassertiefe_2d:standard_name = "sea_floor_depth_below_sea_surface" ;
    Mesh2_face_Gesamtwassertiefe_2d:mesh = "Mesh2" ;
    Mesh2_face_Gesamtwassertiefe_2d:location = "face" ;

// -----------------------------------------------------------------------------
// -----------------------------------------------------------------------------
// -----------------------------------------------------------------------------
// ---------------  Here come non-standart variables... ------------------------
// -----------------------------------------------------------------------------
// -----------------------------------------------------------------------------
// -----------------------------------------------------------------------------

float Mesh2_face_WaveHeight_2d(nMesh2_data_time, nMesh2_face) ;
    Mesh2_face_WaveHeight_2d:long_name = "wave_height, Face (Polygon)" ; 
    Mesh2_face_WaveHeight_2d:units = "m" ; 
    Mesh2_face_WaveHeight_2d:name_id = 840 ; 
    Mesh2_face_WaveHeight_2d:_FillValue = 1.e+31f ; 
    Mesh2_face_WaveHeight_2d:cell_measures = "area: Mesh2_face_wet_area" ; 
    Mesh2_face_WaveHeight_2d:cell_methods = "nMesh2_data_time: point area: mean" ; 
    Mesh2_face_WaveHeight_2d:coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ;
    Mesh2_face_WaveHeight_2d:grid_mapping = "Mesh2_crs" ; 
    Mesh2_face_WaveHeight_2d:standard_name = 'wave_height' ; 
    Mesh2_face_WaveHeight_2d:mesh = "Mesh2" ; 
    Mesh2_face_WaveHeight_2d:location = "face" ;
    // Mesh2_face_WaveHeight_2d:davit_role = "visualization_variable" ;

float Mesh2_face_SedimentFluxAtSoil_2d (nMesh2_data_time, nMesh2_face) ;
    Mesh2_face_SedimentFluxAtSoil_2d: long_name = 'concentration_of_SPM_upward_flux_at_soil_surface, Face (Polygon)' ; 
    Mesh2_face_SedimentFluxAtSoil_2d: standard_name = 'concentration_of_SPM_upward_flux_at_soil_surface' ; 
    Mesh2_face_SedimentFluxAtSoil_2d: units = '???' ;
    // in PHYDEF units: kg/m2/s
    Mesh2_face_SedimentFluxAtSoil_2d: name_id = 1478 ; 
    Mesh2_face_SedimentFluxAtSoil_2d: _FillValue = 1.e+31f ; 
    Mesh2_face_SedimentFluxAtSoil_2d: mesh = "Mesh2" ; 
    Mesh2_face_SedimentFluxAtSoil_2d: location = "face" ;
    // Mesh2_face_SedimentFluxAtSoil_2d: cell_measures = "area: Mesh2_face_wet_area" ; 
    // Mesh2_face_SedimentFluxAtSoil_2d: cell_methods = "nMesh2_data_time: point area: mean" ; 
    Mesh2_face_SedimentFluxAtSoil_2d: coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ;
    Mesh2_face_SedimentFluxAtSoil_2d: grid_mapping = "Mesh2_crs" ; 

float Mesh2_face_RadiactiveFluxAtSurface_2d (nMesh2_data_time, nMesh2_face) ;
    Mesh2_face_RadiactiveFluxAtSurface_2d: long_name = 'surface_downwelling_photosynthetic_radiative_flux, Face (Polygon)' ; 
    Mesh2_face_RadiactiveFluxAtSurface_2d: standard_name = 'surface_downwelling_photosynthetic_radiative_flux' ; 
    Mesh2_face_RadiactiveFluxAtSurface_2d: units = 'W/m**2' ;
    Mesh2_face_RadiactiveFluxAtSurface_2d: name_id = 1153 ; 
    Mesh2_face_RadiactiveFluxAtSurface_2d: _FillValue = 1.e+31f ; 
    Mesh2_face_RadiactiveFluxAtSurface_2d: mesh = "Mesh2" ; 
    Mesh2_face_RadiactiveFluxAtSurface_2d: location = "face" ;
    // Mesh2_face_RadiactiveFluxAtSurface_2d: cell_measures = "area: Mesh2_face_wet_area" ; 
    // Mesh2_face_RadiactiveFluxAtSurface_2d: cell_methods = "nMesh2_data_time: point area: mean" ; 
    Mesh2_face_RadiactiveFluxAtSurface_2d: coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ;
    Mesh2_face_RadiactiveFluxAtSurface_2d: grid_mapping = "Mesh2_crs" ; 

float Mesh2_face_TemperatureAtSoil_2d (nMesh2_data_time, nMesh2_face) ;
    Mesh2_face_TemperatureAtSoil_2d: long_name = 'temperature_at_soil_surface, Face (Polygon)' ; 
    Mesh2_face_TemperatureAtSoil_2d: standard_name = 'temperature_at_soil_surface' ; 
    Mesh2_face_TemperatureAtSoil_2d: units = 'degr.C.' ;
    Mesh2_face_TemperatureAtSoil_2d: name_id = 6 ; 
    Mesh2_face_TemperatureAtSoil_2d: _FillValue = 1.e+31f ; 
    Mesh2_face_TemperatureAtSoil_2d: mesh = "Mesh2" ; 
    Mesh2_face_TemperatureAtSoil_2d: location = "face" ;
    // Mesh2_face_TemperatureAtSoil_2d: cell_measures = "area: Mesh2_face_wet_area" ; 
    // Mesh2_face_TemperatureAtSoil_2d: cell_methods = "nMesh2_data_time: point area: mean" ; 
    Mesh2_face_TemperatureAtSoil_2d: coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ;
    Mesh2_face_TemperatureAtSoil_2d: grid_mapping = "Mesh2_crs" ;

float Mesh2_face_TurbulentMomentumDiffusivityAtSoil_2d (nMesh2_data_time, nMesh2_face) ;
    Mesh2_face_TurbulentMomentumDiffusivityAtSoil_2d: long_name = 'turbulent_diffusivity_of_momentum_at_soil_surface, Face (Polygon)' ; 
    Mesh2_face_TurbulentMomentumDiffusivityAtSoil_2d: standard_name = 'turbulent_diffusivity_of_momentum_at_soil_surface' ; 
    Mesh2_face_TurbulentMomentumDiffusivityAtSoil_2d: units = 'm**2/s' ;
    Mesh2_face_TurbulentMomentumDiffusivityAtSoil_2d: name_id = 873 ; 
    Mesh2_face_TurbulentMomentumDiffusivityAtSoil_2d: _FillValue = 1.e+31f ; 
    Mesh2_face_TurbulentMomentumDiffusivityAtSoil_2d: mesh = "Mesh2" ; 
    Mesh2_face_TurbulentMomentumDiffusivityAtSoil_2d: location = "face" ;
    // Mesh2_face_TurbulentMomentumDiffusivityAtSoil_2d: cell_measures = "area: Mesh2_face_wet_area" ; 
    // Mesh2_face_TurbulentMomentumDiffusivityAtSoil_2d: cell_methods = "nMesh2_data_time: point area: mean" ; 
    Mesh2_face_TurbulentMomentumDiffusivityAtSoil_2d: coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ;
    Mesh2_face_TurbulentMomentumDiffusivityAtSoil_2d: grid_mapping = "Mesh2_crs" ;

float Mesh2_face_WaveSpreadingDirection_2d (nMesh2_data_time, nMesh2_face) ;
    Mesh2_face_WaveSpreadingDirection_2d: long_name = 'wave_direction, Face (Polygon)' ; 
    Mesh2_face_WaveSpreadingDirection_2d: standard_name = 'wave_direction' ; 
    Mesh2_face_WaveSpreadingDirection_2d: units = 'rad' ;
    // in PHYDEF units = 'degree'
    Mesh2_face_WaveSpreadingDirection_2d: name_id = 1005 ; 
    Mesh2_face_WaveSpreadingDirection_2d: _FillValue = 1.e+31f ; 
    Mesh2_face_WaveSpreadingDirection_2d: mesh = "Mesh2" ; 
    Mesh2_face_WaveSpreadingDirection_2d: location = "face" ;
    // Mesh2_face_WaveSpreadingDirection_2d: cell_measures = "area: Mesh2_face_wet_area" ; 
    // Mesh2_face_WaveSpreadingDirection_2d: cell_methods = "nMesh2_data_time: point area: mean" ; 
    Mesh2_face_WaveSpreadingDirection_2d: coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ;
    Mesh2_face_WaveSpreadingDirection_2d: grid_mapping = "Mesh2_crs" ;

float Mesh2_face_WaveNumber_2d (nMesh2_data_time, nMesh2_face) ;
    Mesh2_face_WaveNumber_2d: long_name = 'wave_number, Face (Polygon)' ; 
    Mesh2_face_WaveNumber_2d: standard_name = 'wave_number' ; 
    Mesh2_face_WaveNumber_2d: units = '1/m' ;
    // in PHYDEF units = 'rad/m'
    Mesh2_face_WaveNumber_2d: name_id = 845 ; 
    Mesh2_face_WaveNumber_2d: _FillValue = 1.e+31f ; 
    Mesh2_face_WaveNumber_2d: mesh = "Mesh2" ; 
    Mesh2_face_WaveNumber_2d: location = "face" ;
    // Mesh2_face_WaveNumber_2d: cell_measures = "area: Mesh2_face_wet_area" ; 
    // Mesh2_face_WaveNumber_2d: cell_methods = "nMesh2_data_time: point area: mean" ; 
    Mesh2_face_WaveNumber_2d: coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ;
    Mesh2_face_WaveNumber_2d: grid_mapping = "Mesh2_crs" ;

float Mesh2_face_MeanWavePeriod_2d (nMesh2_data_time, nMesh2_face) ;
    Mesh2_face_MeanWavePeriod_2d: long_name = 'wave_period, Face (Polygon)' ; 
    Mesh2_face_MeanWavePeriod_2d: standard_name = 'wave_period' ; 
    Mesh2_face_MeanWavePeriod_2d: units = 's' ;
    Mesh2_face_MeanWavePeriod_2d: name_id = 1000 ; 
    Mesh2_face_MeanWavePeriod_2d: _FillValue = 1.e+31f ; 
    Mesh2_face_MeanWavePeriod_2d: mesh = "Mesh2" ; 
    Mesh2_face_MeanWavePeriod_2d: location = "face" ;
    // Mesh2_face_MeanWavePeriod_2d: cell_measures = "area: Mesh2_face_wet_area" ; 
    // Mesh2_face_MeanWavePeriod_2d: cell_methods = "nMesh2_data_time: point area: mean" ; 
    Mesh2_face_MeanWavePeriod_2d: coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ;
    Mesh2_face_MeanWavePeriod_2d: grid_mapping = "Mesh2_crs" ;

float Mesh2_face_WindVelocityAt10m_x_2d(nMesh2_data_time, nMesh2_face) ;
    Mesh2_face_WindVelocityAt10m_x_2d: long_name = "wind_velocityAt10m (x-Komponente), Face (Polygon)" ; 
    Mesh2_face_WindVelocityAt10m_x_2d: units = "m s-1" ; 
    Mesh2_face_WindVelocityAt10m_x_2d: name_id = 557 ; 
    Mesh2_face_WindVelocityAt10m_x_2d: _FillValue = 1.e+31f ; 
    Mesh2_face_WindVelocityAt10m_x_2d: cell_methods = "nMesh2_data_time: point nMesh2_layer_2d: mean area: point" ; 
    Mesh2_face_WindVelocityAt10m_x_2d: coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ; 
    Mesh2_face_WindVelocityAt10m_x_2d: grid_mapping = "Mesh2_crs" ; 
    Mesh2_face_WindVelocityAt10m_x_2d: standard_name = "wind_x_velocityAt10m" ; 
    Mesh2_face_WindVelocityAt10m_x_2d: mesh = "Mesh2" ; 
    Mesh2_face_WindVelocityAt10m_x_2d: location = "face" ; 
    // Mesh2_face_WindVelocityAt10m_x_2d :davit_role = "visualization_variable" ;

float Mesh2_face_WindVelocityAt10m_y_2d(nMesh2_data_time, nMesh2_face) ;
    Mesh2_face_WindVelocityAt10m_y_2d: long_name = "wind_velocityAt10m (y-Komponente), Face (Polygon)" ; 
    Mesh2_face_WindVelocityAt10m_y_2d: units = "m s-1" ; 
    Mesh2_face_WindVelocityAt10m_y_2d: name_id = 558 ; 
    Mesh2_face_WindVelocityAt10m_y_2d: _FillValue = 1.e+31f ; 
    Mesh2_face_WindVelocityAt10m_y_2d: cell_methods = "nMesh2_data_time: point nMesh2_layer_2d: mean area: point" ; 
    Mesh2_face_WindVelocityAt10m_y_2d: coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ; 
    Mesh2_face_WindVelocityAt10m_y_2d: grid_mapping = "Mesh2_crs" ; 
    Mesh2_face_WindVelocityAt10m_y_2d: standard_name = "wind_y_velocityAt10m" ; 
    Mesh2_face_WindVelocityAt10m_y_2d: mesh = "Mesh2" ; 
    Mesh2_face_WindVelocityAt10m_y_2d: location = "face" ; 
    // Mesh2_face_WindVelocityAt10m_y_2d: davit_role = "visualization_variable" ;

float Mesh2_face_WindVelocityAt10m_m_2d(nMesh2_data_time, nMesh2_face) ;
    Mesh2_face_WindVelocityAt10m_m_2d: long_name = "wind_velocityAt10m (Betrag), Face (Polygon)" ; 
    Mesh2_face_WindVelocityAt10m_m_2d: units = "m s-1" ; 
    Mesh2_face_WindVelocityAt10m_m_2d: name_id = 906 ; 
    Mesh2_face_WindVelocityAt10m_m_2d: _FillValue = 1.e+31f ; 
    Mesh2_face_WindVelocityAt10m_m_2d: cell_methods = "nMesh2_data_time: point nMesh2_layer_2d: mean area: point" ; 
    Mesh2_face_WindVelocityAt10m_m_2d: coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ; 
    Mesh2_face_WindVelocityAt10m_m_2d: grid_mapping = "Mesh2_crs" ; 
    Mesh2_face_WindVelocityAt10m_m_2d: standard_name = "magnitude_of_wind_velocityAt10m" ; 
    Mesh2_face_WindVelocityAt10m_m_2d: mesh = "Mesh2" ; 
    Mesh2_face_WindVelocityAt10m_m_2d: location = "face" ; 
    // Mesh2_face_WindVelocityAt10m_m_2d: davit_role = "visualization_variable" ;

float Mesh2_face_WaterVelocityAtSoil_x_2d(nMesh2_data_time, nMesh2_face) ;
    Mesh2_face_WaterVelocityAtSoil_x_2d: long_name = "velocityAtSoil_surface (x-Komponente), Face (Polygon)" ; 
    Mesh2_face_WaterVelocityAtSoil_x_2d: units = "m s-1" ; 
    Mesh2_face_WaterVelocityAtSoil_x_2d: name_id = 14 ; 
    Mesh2_face_WaterVelocityAtSoil_x_2d: _FillValue = 1.e+31f ; 
    Mesh2_face_WaterVelocityAtSoil_x_2d: cell_methods = "nMesh2_data_time: point nMesh2_layer_2d: mean area: point" ; 
    Mesh2_face_WaterVelocityAtSoil_x_2d: coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ; 
    Mesh2_face_WaterVelocityAtSoil_x_2d: grid_mapping = "Mesh2_crs" ; 
    Mesh2_face_WaterVelocityAtSoil_x_2d: standard_name = "x_velocityAtSoil_surface" ; 
    Mesh2_face_WaterVelocityAtSoil_x_2d: mesh = "Mesh2" ; 
    Mesh2_face_WaterVelocityAtSoil_x_2d: location = "face" ; 
    // Mesh2_face_WaterVelocityAtSoil_x_2d :davit_role = "visualization_variable" ;

float Mesh2_face_WaterVelocityAtSoil_y_2d(nMesh2_data_time, nMesh2_face) ;
    Mesh2_face_WaterVelocityAtSoil_y_2d: long_name = "velocityAtSoil_surface (y-Komponente), Face (Polygon)" ; 
    Mesh2_face_WaterVelocityAtSoil_y_2d: units = "m s-1" ; 
    Mesh2_face_WaterVelocityAtSoil_y_2d: name_id = 15 ; 
    Mesh2_face_WaterVelocityAtSoil_y_2d: _FillValue = 1.e+31f ; 
    Mesh2_face_WaterVelocityAtSoil_y_2d: cell_methods = "nMesh2_data_time: point nMesh2_layer_2d: mean area: point" ; 
    Mesh2_face_WaterVelocityAtSoil_y_2d: coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ; 
    Mesh2_face_WaterVelocityAtSoil_y_2d: grid_mapping = "Mesh2_crs" ; 
    Mesh2_face_WaterVelocityAtSoil_y_2d: standard_name = "y_velocityAtSoil_surface" ; 
    Mesh2_face_WaterVelocityAtSoil_y_2d: mesh = "Mesh2" ; 
    Mesh2_face_WaterVelocityAtSoil_y_2d: location = "face" ; 
    // Mesh2_face_WaterVelocityAtSoil_y_2d: davit_role = "visualization_variable" ;

float Mesh2_face_WaterVelocityAtSoil_m_2d(nMesh2_data_time, nMesh2_face) ;
    Mesh2_face_WaterVelocityAtSoil_m_2d: long_name = "velocityAtSoil_surface (Betrag), Face (Polygon)" ; 
    Mesh2_face_WaterVelocityAtSoil_m_2d: units = "m s-1" ; 
    Mesh2_face_WaterVelocityAtSoil_m_2d: name_id = 2 ; 
    Mesh2_face_WaterVelocityAtSoil_m_2d: _FillValue = 1.e+31f ; 
    Mesh2_face_WaterVelocityAtSoil_m_2d: cell_methods = "nMesh2_data_time: point nMesh2_layer_2d: mean area: point" ; 
    Mesh2_face_WaterVelocityAtSoil_m_2d: coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ; 
    Mesh2_face_WaterVelocityAtSoil_m_2d: grid_mapping = "Mesh2_crs" ; 
    Mesh2_face_WaterVelocityAtSoil_m_2d: standard_name = "magnitude_of_velocityAtSoil_surface" ; 
    Mesh2_face_WaterVelocityAtSoil_m_2d: mesh = "Mesh2" ; 
    Mesh2_face_WaterVelocityAtSoil_m_2d: location = "face" ; 
    // Mesh2_face_WaterVelocityAtSoil_m_2d: davit_role = "visualization_variable" ;