netcdf nsbs_davit {
dimensions:
	nMesh2_node = 10918 ;
	nMesh2_edge = 20998 ;
	nMesh2_face = 10061 ;
	nMaxMesh2_face_nodes = 4 ;
	two = 2 ;
	three = 3 ;
	nMesh2_time = 1 ;
	nMesh2_data_time = UNLIMITED ; // (5 currently)
	nMesh2_layer_2d = 1 ;
	nMesh2_layer_3d = 30 ;
	nMesh2_class_names_strlen = 20 ;
	nMesh2_suspension_classes = 1 ;
variables:
	int Mesh2_crs ;
		Mesh2_crs:epsg_code = "EPSG:4326" ;
		Mesh2_crs:comment = "LON, LAT : WGS84, EPSG:4326" ;
		Mesh2_crs:grid_mapping_name = "latitude_longitude" ;
		Mesh2_crs:longitude_of_prime_meridian = 0. ;
		Mesh2_crs:semi_major_axis = 6378137. ;
		Mesh2_crs:inverse_flattening = 298.257223563 ;
	double Mesh2_node_lon(nMesh2_node) ;
		Mesh2_node_lon:long_name = "geografische Laenge der 2D-Gitter-Knoten" ;
		Mesh2_node_lon:units = "degrees_east" ;
		Mesh2_node_lon:name_id = 1653 ;
		Mesh2_node_lon:standard_name = "longitude" ;
	double Mesh2_node_lat(nMesh2_node) ;
		Mesh2_node_lat:long_name = "geografische Breite der 2D-Gitter-Knoten" ;
		Mesh2_node_lat:units = "degrees_north" ;
		Mesh2_node_lat:name_id = 1652 ;
		Mesh2_node_lat:standard_name = "latitude" ;
	double Mesh2_edge_lon(nMesh2_edge) ;
		Mesh2_edge_lon:long_name = "geografische Laenge der 2D-Gitter-Kanten, Kantenmitte" ;
		Mesh2_edge_lon:units = "degrees_east" ;
		Mesh2_edge_lon:name_id = 1653 ;
		Mesh2_edge_lon:bounds = "Mesh2_edge_lon_bnd" ;
		Mesh2_edge_lon:standard_name = "longitude" ;
	double Mesh2_edge_lat(nMesh2_edge) ;
		Mesh2_edge_lat:long_name = "geografische Breite der 2D-Gitter-Kanten, Kantenmitte" ;
		Mesh2_edge_lat:units = "degrees_north" ;
		Mesh2_edge_lat:name_id = 1652 ;
		Mesh2_edge_lat:bounds = "Mesh2_edge_lat_bnd" ;
		Mesh2_edge_lat:standard_name = "latitude" ;
	double Mesh2_face_lon(nMesh2_face) ;
		Mesh2_face_lon:long_name = "geografische Laenge der 2D-Gitter-Faces (Polygone), Schwerpunkt" ;
		Mesh2_face_lon:units = "degrees_east" ;
		Mesh2_face_lon:name_id = 1653 ;
		Mesh2_face_lon:bounds = "Mesh2_face_lon_bnd" ;
		Mesh2_face_lon:standard_name = "longitude" ;
	double Mesh2_face_lat(nMesh2_face) ;
		Mesh2_face_lat:long_name = "geografische Breite der 2D-Gitter-Faces (Polygone), Schwerpunkt" ;
		Mesh2_face_lat:units = "degrees_north" ;
		Mesh2_face_lat:name_id = 1652 ;
		Mesh2_face_lat:bounds = "Mesh2_face_lat_bnd" ;
		Mesh2_face_lat:standard_name = "latitude" ;
	double Mesh2_face_center_lon(nMesh2_face) ;
		Mesh2_face_center_lon:long_name = "geografische Laenge der 2D-Gitter-Faces (Polygone), Umkreismittelpunkt" ;
		Mesh2_face_center_lon:units = "degrees_east" ;
		Mesh2_face_center_lon:name_id = 1653 ;
		Mesh2_face_center_lon:standard_name = "longitude" ;
	double Mesh2_face_center_lat(nMesh2_face) ;
		Mesh2_face_center_lat:long_name = "geografische Breite der 2D-Gitter-faces (Polygone), Umkreismittelpunkt" ;
		Mesh2_face_center_lat:units = "degrees_north" ;
		Mesh2_face_center_lat:name_id = 1652 ;
		Mesh2_face_center_lat:standard_name = "latitude" ;
	double Mesh2_edge_lon_bnd(nMesh2_edge, two) ;
	double Mesh2_edge_lat_bnd(nMesh2_edge, two) ;
	double Mesh2_face_lon_bnd(nMesh2_face, nMaxMesh2_face_nodes) ;
		Mesh2_face_lon_bnd:_FillValue = -999. ;
	double Mesh2_face_lat_bnd(nMesh2_face, nMaxMesh2_face_nodes) ;
		Mesh2_face_lat_bnd:_FillValue = -999. ;
	int Mesh2 ;
		Mesh2:long_name = "UnTRIM Gitternetz, Vierecke, kein SubGrid" ;
		Mesh2:cf_role = "mesh_topology" ;
		Mesh2:dimensionality = 2 ;
		Mesh2:node_coordinates = "Mesh2_node_lon Mesh2_node_lat Mesh2_node_x Mesh2_node_y" ;
		Mesh2:edge_coordinates = "Mesh2_edge_lon Mesh2_edge_lat Mesh2_edge_x Mesh2_edge_y" ;
		Mesh2:face_coordinates = "Mesh2_face_lon Mesh2_face_lat Mesh2_face_x Mesh2_face_y Mesh2_face_center_lon Mesh2_face_center_lat Mesh2_face_center_x Mesh2_face_center_y " ;
		Mesh2:edge_node_connectivity = "Mesh2_edge_nodes" ;
		Mesh2:edge_face_connectivity = "Mesh2_edge_faces" ;
		Mesh2:face_node_connectivity = "Mesh2_face_nodes" ;
		Mesh2:face_edge_connectivity = "Mesh2_face_edges" ;
	int Mesh2_edge_nodes(nMesh2_edge, two) ;
		Mesh2_edge_nodes:long_name = "Knotenverzeichnis der Kanten, Anfangs- und Endpunkt" ;
		Mesh2_edge_nodes:cf_role = "edge_node_connectivity" ;
		Mesh2_edge_nodes:start_index = 0 ;
	int Mesh2_edge_faces(nMesh2_edge, two) ;
		Mesh2_edge_faces:_FillValue = -999 ;
		Mesh2_edge_faces:long_name = "Face- (Polygon-) Verzeichnis der Kanten, linker und rechter Nachbar" ;
		Mesh2_edge_faces:cf_role = "edge_face_connectivity" ;
		Mesh2_edge_faces:start_index = 0 ;
	int Mesh2_face_nodes(nMesh2_face, nMaxMesh2_face_nodes) ;
		Mesh2_face_nodes:_FillValue = -999 ;
		Mesh2_face_nodes:long_name = "Knotenverzeichnis der Faces (Polygone),entgegen dem Uhrzeigersinn" ;
		Mesh2_face_nodes:cf_role = "face_node_connectivity" ;
		Mesh2_face_nodes:start_index = 0 ;
	int Mesh2_face_edges(nMesh2_face, nMaxMesh2_face_nodes) ;
		Mesh2_face_edges:_FillValue = -999 ;
		Mesh2_face_edges:long_name = "Kantenverzeichnis der Faces (Polygone),entgegen dem Uhrzeigersinn" ;
		Mesh2_face_edges:cf_role = "face_edge_connectivity" ;
		Mesh2_face_edges:start_index = 0 ;
	double nMesh2_time(nMesh2_time) ;
		nMesh2_time:bounds = "nMesh2_time_bnd" ;
		nMesh2_time:long_name = "time" ;
		nMesh2_time:standard_name = "time" ;
		nMesh2_time:name_id = 1640 ;
		nMesh2_time:units = "seconds since 2008-01-02 00:00:00 01:00" ;
		nMesh2_time:calendar = "gregorian" ;
		nMesh2_time:axis = "T" ;
	double nMesh2_time_bnd(nMesh2_time, two) ;
	double nMesh2_data_time(nMesh2_data_time) ;
		nMesh2_data_time:long_name = "time" ;
		nMesh2_data_time:standard_name = "time" ;
		nMesh2_data_time:name_id = 1640 ;
		nMesh2_data_time:units = "hours since 2009-01-02 00:00:00 01:00" ;
		nMesh2_data_time:calendar = "gregorian" ;
		nMesh2_data_time:axis = "T" ;
	float Mesh2_face_z_face_3d(nMesh2_data_time, nMesh2_layer_3d, nMesh2_face) ;
		Mesh2_face_z_face_3d:positive = "down" ;
		Mesh2_face_z_face_3d:bounds = "Mesh2_face_z_face_bnd_3d" ;
		Mesh2_face_z_face_3d:long_name = "z_face [ face ]" ;
		Mesh2_face_z_face_3d:standard_name = "depth" ;
		Mesh2_face_z_face_3d:name_id = 1702 ;
		Mesh2_face_z_face_3d:units = "m" ;
	float Mesh2_face_z_face_bnd_3d(nMesh2_data_time, nMesh2_layer_3d, nMesh2_face, two) ;
		Mesh2_face_z_face_bnd_3d:name_id = 1703 ;
	float Mesh2_edge_z_edge_3d(nMesh2_data_time, nMesh2_layer_3d, nMesh2_edge) ;
		Mesh2_edge_z_edge_3d:positive = "down" ;
		Mesh2_edge_z_edge_3d:bounds = "Mesh2_edge_z_edge_bnd_3d" ;
		Mesh2_edge_z_edge_3d:long_name = "z_edge [ edge ]" ;
		Mesh2_edge_z_edge_3d:standard_name = "depth" ;
		Mesh2_edge_z_edge_3d:name_id = 1707 ;
		Mesh2_edge_z_edge_3d:units = "m" ;
	float Mesh2_edge_z_edge_bnd_3d(nMesh2_data_time, nMesh2_layer_3d, nMesh2_edge, two) ;
		Mesh2_edge_z_edge_bnd_3d:name_id = 1708 ;
	float Mesh2_face_RadiactiveFluxAtSurface_2d(nMesh2_data_time, nMesh2_face) ;
		Mesh2_face_RadiactiveFluxAtSurface_2d:_FillValue = 1.e+31f ;
		Mesh2_face_RadiactiveFluxAtSurface_2d:grid_mapping = "Mesh2_crs" ;
		Mesh2_face_RadiactiveFluxAtSurface_2d:coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ;
		Mesh2_face_RadiactiveFluxAtSurface_2d:long_name = "surface_downwelling_photosynthetic_radiative_flux, Face (Polygon)" ;
		Mesh2_face_RadiactiveFluxAtSurface_2d:standard_name = "surface_downwelling_photosynthetic_radiative_flux" ;
		Mesh2_face_RadiactiveFluxAtSurface_2d:mesh = "Mesh2" ;
		Mesh2_face_RadiactiveFluxAtSurface_2d:name_id = 1153 ;
		Mesh2_face_RadiactiveFluxAtSurface_2d:location = "face" ;
		Mesh2_face_RadiactiveFluxAtSurface_2d:units = "W/m**2" ;
	double Mesh2_face_depth_2d(nMesh2_time, nMesh2_face) ;
		Mesh2_face_depth_2d:_FillValue = 1.e+31 ;
		Mesh2_face_depth_2d:grid_mapping = "Mesh2_crs" ;
		Mesh2_face_depth_2d:coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ;
		Mesh2_face_depth_2d:valid_range = -8848., 11034. ;
		Mesh2_face_depth_2d:long_name = "Topographie" ;
		Mesh2_face_depth_2d:standard_name = "sea_floor_depth_below_geoid" ;
		Mesh2_face_depth_2d:mesh = "Mesh2" ;
		Mesh2_face_depth_2d:name_id = 17 ;
		Mesh2_face_depth_2d:location = "face" ;
		Mesh2_face_depth_2d:cell_methods = "nMesh2_time: mean area: mean" ;
		Mesh2_face_depth_2d:units = "m" ;
		Mesh2_face_depth_2d:cell_measures = "area: Mesh2_face_area" ;
	float Mesh2_face_WaveNumber_2d(nMesh2_data_time, nMesh2_face) ;
		Mesh2_face_WaveNumber_2d:_FillValue = 1.e+31f ;
		Mesh2_face_WaveNumber_2d:grid_mapping = "Mesh2_crs" ;
		Mesh2_face_WaveNumber_2d:coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ;
		Mesh2_face_WaveNumber_2d:long_name = "wave_number, Face (Polygon)" ;
		Mesh2_face_WaveNumber_2d:standard_name = "wave_number" ;
		Mesh2_face_WaveNumber_2d:mesh = "Mesh2" ;
		Mesh2_face_WaveNumber_2d:name_id = 845 ;
		Mesh2_face_WaveNumber_2d:location = "face" ;
		Mesh2_face_WaveNumber_2d:units = "1/m" ;
	float Mesh2_face_Stroemungsgeschwindigkeit_x_2d(nMesh2_data_time, nMesh2_layer_2d, nMesh2_face) ;
		Mesh2_face_Stroemungsgeschwindigkeit_x_2d:_FillValue = 1.e+31f ;
		Mesh2_face_Stroemungsgeschwindigkeit_x_2d:grid_mapping = "Mesh2_crs" ;
		Mesh2_face_Stroemungsgeschwindigkeit_x_2d:coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat Mesh2_face_z_face_2d" ;
		Mesh2_face_Stroemungsgeschwindigkeit_x_2d:long_name = "Stroemungsgeschwindigkeit (x-Komponente), Face (Polygon)" ;
		Mesh2_face_Stroemungsgeschwindigkeit_x_2d:standard_name = "sea_water_x_velocity" ;
		Mesh2_face_Stroemungsgeschwindigkeit_x_2d:cell_methods = "nMesh2_data_time: point nMesh2_layer_2d: mean area: point" ;
		Mesh2_face_Stroemungsgeschwindigkeit_x_2d:name_id = 2 ;
		Mesh2_face_Stroemungsgeschwindigkeit_x_2d:location = "face" ;
		Mesh2_face_Stroemungsgeschwindigkeit_x_2d:units = "m s-1" ;
		Mesh2_face_Stroemungsgeschwindigkeit_x_2d:mesh = "Mesh2" ;
	float Mesh2_face_WaveHeight_2d(nMesh2_data_time, nMesh2_face) ;
		Mesh2_face_WaveHeight_2d:_FillValue = 1.e+31f ;
		Mesh2_face_WaveHeight_2d:grid_mapping = "Mesh2_crs" ;
		Mesh2_face_WaveHeight_2d:cell_measures = "area: Mesh2_face_wet_area" ;
		Mesh2_face_WaveHeight_2d:coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ;
		Mesh2_face_WaveHeight_2d:long_name = "wave_height, Face (Polygon)" ;
		Mesh2_face_WaveHeight_2d:standard_name = "wave_height" ;
		Mesh2_face_WaveHeight_2d:cell_methods = "nMesh2_data_time: point area: mean" ;
		Mesh2_face_WaveHeight_2d:name_id = 840 ;
		Mesh2_face_WaveHeight_2d:location = "face" ;
		Mesh2_face_WaveHeight_2d:units = "m" ;
		Mesh2_face_WaveHeight_2d:mesh = "Mesh2" ;
	float Mesh2_face_SedimentFluxAtSoil_2d(nMesh2_data_time, nMesh2_face) ;
		Mesh2_face_SedimentFluxAtSoil_2d:_FillValue = 1.e+31f ;
		Mesh2_face_SedimentFluxAtSoil_2d:grid_mapping = "Mesh2_crs" ;
		Mesh2_face_SedimentFluxAtSoil_2d:coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ;
		Mesh2_face_SedimentFluxAtSoil_2d:long_name = "concentration_of_SPM_upward_flux_at_soil_surface, Face (Polygon)" ;
		Mesh2_face_SedimentFluxAtSoil_2d:standard_name = "concentration_of_SPM_upward_flux_at_soil_surface" ;
		Mesh2_face_SedimentFluxAtSoil_2d:mesh = "Mesh2" ;
		Mesh2_face_SedimentFluxAtSoil_2d:name_id = 1478 ;
		Mesh2_face_SedimentFluxAtSoil_2d:location = "face" ;
		Mesh2_face_SedimentFluxAtSoil_2d:units = "???" ;
	float Mesh2_face_TurbulentMomentumDiffusivityAtSoil_2d(nMesh2_data_time, nMesh2_face) ;
		Mesh2_face_TurbulentMomentumDiffusivityAtSoil_2d:_FillValue = 1.e+31f ;
		Mesh2_face_TurbulentMomentumDiffusivityAtSoil_2d:grid_mapping = "Mesh2_crs" ;
		Mesh2_face_TurbulentMomentumDiffusivityAtSoil_2d:coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ;
		Mesh2_face_TurbulentMomentumDiffusivityAtSoil_2d:long_name = "turbulent_diffusivity_of_momentum_at_soil_surface, Face (Polygon)" ;
		Mesh2_face_TurbulentMomentumDiffusivityAtSoil_2d:standard_name = "turbulent_diffusivity_of_momentum_at_soil_surface" ;
		Mesh2_face_TurbulentMomentumDiffusivityAtSoil_2d:mesh = "Mesh2" ;
		Mesh2_face_TurbulentMomentumDiffusivityAtSoil_2d:name_id = 873 ;
		Mesh2_face_TurbulentMomentumDiffusivityAtSoil_2d:location = "face" ;
		Mesh2_face_TurbulentMomentumDiffusivityAtSoil_2d:units = "m**2/s" ;
	float Mesh2_face_TemperatureAtSoil_2d(nMesh2_data_time, nMesh2_face) ;
		Mesh2_face_TemperatureAtSoil_2d:_FillValue = 1.e+31f ;
		Mesh2_face_TemperatureAtSoil_2d:grid_mapping = "Mesh2_crs" ;
		Mesh2_face_TemperatureAtSoil_2d:coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ;
		Mesh2_face_TemperatureAtSoil_2d:long_name = "temperature_at_soil_surface, Face (Polygon)" ;
		Mesh2_face_TemperatureAtSoil_2d:standard_name = "temperature_at_soil_surface" ;
		Mesh2_face_TemperatureAtSoil_2d:mesh = "Mesh2" ;
		Mesh2_face_TemperatureAtSoil_2d:name_id = 6 ;
		Mesh2_face_TemperatureAtSoil_2d:location = "face" ;
		Mesh2_face_TemperatureAtSoil_2d:units = "degr.C." ;
	float Mesh2_face_WaterVelocityAtSoil_y_2d(nMesh2_data_time, nMesh2_face) ;
		Mesh2_face_WaterVelocityAtSoil_y_2d:_FillValue = 1.e+31f ;
		Mesh2_face_WaterVelocityAtSoil_y_2d:grid_mapping = "Mesh2_crs" ;
		Mesh2_face_WaterVelocityAtSoil_y_2d:coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ;
		Mesh2_face_WaterVelocityAtSoil_y_2d:long_name = "velocityAtSoil_surface (y-Komponente), Face (Polygon)" ;
		Mesh2_face_WaterVelocityAtSoil_y_2d:standard_name = "y_velocityAtSoil_surface" ;
		Mesh2_face_WaterVelocityAtSoil_y_2d:cell_methods = "nMesh2_data_time: point nMesh2_layer_2d: mean area: point" ;
		Mesh2_face_WaterVelocityAtSoil_y_2d:name_id = 15 ;
		Mesh2_face_WaterVelocityAtSoil_y_2d:location = "face" ;
		Mesh2_face_WaterVelocityAtSoil_y_2d:units = "m s-1" ;
		Mesh2_face_WaterVelocityAtSoil_y_2d:mesh = "Mesh2" ;
	float Mesh2_face_WaveSpreadingDirection_2d(nMesh2_data_time, nMesh2_face) ;
		Mesh2_face_WaveSpreadingDirection_2d:_FillValue = 1.e+31f ;
		Mesh2_face_WaveSpreadingDirection_2d:grid_mapping = "Mesh2_crs" ;
		Mesh2_face_WaveSpreadingDirection_2d:coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ;
		Mesh2_face_WaveSpreadingDirection_2d:long_name = "wave_direction, Face (Polygon)" ;
		Mesh2_face_WaveSpreadingDirection_2d:standard_name = "wave_direction" ;
		Mesh2_face_WaveSpreadingDirection_2d:mesh = "Mesh2" ;
		Mesh2_face_WaveSpreadingDirection_2d:name_id = 1005 ;
		Mesh2_face_WaveSpreadingDirection_2d:location = "face" ;
		Mesh2_face_WaveSpreadingDirection_2d:units = "rad" ;
	float Mesh2_face_MeanWavePeriod_2d(nMesh2_data_time, nMesh2_face) ;
		Mesh2_face_MeanWavePeriod_2d:_FillValue = 1.e+31f ;
		Mesh2_face_MeanWavePeriod_2d:grid_mapping = "Mesh2_crs" ;
		Mesh2_face_MeanWavePeriod_2d:coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ;
		Mesh2_face_MeanWavePeriod_2d:long_name = "wave_period, Face (Polygon)" ;
		Mesh2_face_MeanWavePeriod_2d:standard_name = "wave_period" ;
		Mesh2_face_MeanWavePeriod_2d:mesh = "Mesh2" ;
		Mesh2_face_MeanWavePeriod_2d:name_id = 1000 ;
		Mesh2_face_MeanWavePeriod_2d:location = "face" ;
		Mesh2_face_MeanWavePeriod_2d:units = "s" ;
	float Mesh2_face_Gesamtwassertiefe_2d(nMesh2_data_time, nMesh2_face) ;
		Mesh2_face_Gesamtwassertiefe_2d:_FillValue = 1.e+31f ;
		Mesh2_face_Gesamtwassertiefe_2d:grid_mapping = "Mesh2_crs" ;
		Mesh2_face_Gesamtwassertiefe_2d:coordinates = "Mesh2_face_lon Mesh2_face_lat Mesh2_face_x Mesh2_face_y" ;
		Mesh2_face_Gesamtwassertiefe_2d:long_name = "Gesamtwassertiefe [ face ]" ;
		Mesh2_face_Gesamtwassertiefe_2d:standard_name = "sea_floor_depth_below_sea_surface" ;
		Mesh2_face_Gesamtwassertiefe_2d:cell_methods = "nMesh2_data_time: point nMesh2_face: mean" ;
		Mesh2_face_Gesamtwassertiefe_2d:name_id = 16 ;
		Mesh2_face_Gesamtwassertiefe_2d:location = "face" ;
		Mesh2_face_Gesamtwassertiefe_2d:units = "m" ;
		Mesh2_face_Gesamtwassertiefe_2d:mesh = "Mesh2" ;
	float Mesh2_face_Temperatur_3d(nMesh2_data_time, nMesh2_layer_3d, nMesh2_face) ;
		Mesh2_face_Temperatur_3d:_FillValue = 1.e+31f ;
		Mesh2_face_Temperatur_3d:grid_mapping = "Mesh2_crs" ;
		Mesh2_face_Temperatur_3d:cell_measures = "area: Mesh2_face_wet_area" ;
		Mesh2_face_Temperatur_3d:coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat Mesh2_face_z_face_3d" ;
		Mesh2_face_Temperatur_3d:long_name = "Temperatur, Face (Polygon)" ;
		Mesh2_face_Temperatur_3d:standard_name = "temperature" ;
		Mesh2_face_Temperatur_3d:cell_methods = "nMesh2_data_time: point nMesh2_layer_3d: mean area: point" ;
		Mesh2_face_Temperatur_3d:name_id = 6 ;
		Mesh2_face_Temperatur_3d:location = "face" ;
		Mesh2_face_Temperatur_3d:units = "degC" ;
		Mesh2_face_Temperatur_3d:mesh = "Mesh2" ;
	float Mesh2_face_WaterVelocityAtSoil_x_2d(nMesh2_data_time, nMesh2_face) ;
		Mesh2_face_WaterVelocityAtSoil_x_2d:_FillValue = 1.e+31f ;
		Mesh2_face_WaterVelocityAtSoil_x_2d:grid_mapping = "Mesh2_crs" ;
		Mesh2_face_WaterVelocityAtSoil_x_2d:coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ;
		Mesh2_face_WaterVelocityAtSoil_x_2d:long_name = "velocityAtSoil_surface (x-Komponente), Face (Polygon)" ;
		Mesh2_face_WaterVelocityAtSoil_x_2d:standard_name = "x_velocityAtSoil_surface" ;
		Mesh2_face_WaterVelocityAtSoil_x_2d:cell_methods = "nMesh2_data_time: point nMesh2_layer_2d: mean area: point" ;
		Mesh2_face_WaterVelocityAtSoil_x_2d:name_id = 14 ;
		Mesh2_face_WaterVelocityAtSoil_x_2d:location = "face" ;
		Mesh2_face_WaterVelocityAtSoil_x_2d:units = "m s-1" ;
		Mesh2_face_WaterVelocityAtSoil_x_2d:mesh = "Mesh2" ;
	float Mesh2_face_Stroemungsgeschwindigkeit_y_2d(nMesh2_data_time, nMesh2_layer_2d, nMesh2_face) ;
		Mesh2_face_Stroemungsgeschwindigkeit_y_2d:_FillValue = 1.e+31f ;
		Mesh2_face_Stroemungsgeschwindigkeit_y_2d:grid_mapping = "Mesh2_crs" ;
		Mesh2_face_Stroemungsgeschwindigkeit_y_2d:coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat Mesh2_face_z_face_2d" ;
		Mesh2_face_Stroemungsgeschwindigkeit_y_2d:long_name = "Stroemungsgeschwindigkeit (y-Komponente), Face (Polygon)" ;
		Mesh2_face_Stroemungsgeschwindigkeit_y_2d:standard_name = "sea_water_y_velocity" ;
		Mesh2_face_Stroemungsgeschwindigkeit_y_2d:cell_methods = "nMesh2_data_time: point nMesh2_layer_2d: mean area: point" ;
		Mesh2_face_Stroemungsgeschwindigkeit_y_2d:name_id = 2 ;
		Mesh2_face_Stroemungsgeschwindigkeit_y_2d:location = "face" ;
		Mesh2_face_Stroemungsgeschwindigkeit_y_2d:units = "m s-1" ;
		Mesh2_face_Stroemungsgeschwindigkeit_y_2d:mesh = "Mesh2" ;
	float Mesh2_face_WindVelocityAt10m_y_2d(nMesh2_data_time, nMesh2_face) ;
		Mesh2_face_WindVelocityAt10m_y_2d:_FillValue = 1.e+31f ;
		Mesh2_face_WindVelocityAt10m_y_2d:grid_mapping = "Mesh2_crs" ;
		Mesh2_face_WindVelocityAt10m_y_2d:coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ;
		Mesh2_face_WindVelocityAt10m_y_2d:long_name = "wind_velocityAt10m (y-Komponente), Face (Polygon)" ;
		Mesh2_face_WindVelocityAt10m_y_2d:standard_name = "wind_y_velocityAt10m" ;
		Mesh2_face_WindVelocityAt10m_y_2d:cell_methods = "nMesh2_data_time: point nMesh2_layer_2d: mean area: point" ;
		Mesh2_face_WindVelocityAt10m_y_2d:name_id = 558 ;
		Mesh2_face_WindVelocityAt10m_y_2d:location = "face" ;
		Mesh2_face_WindVelocityAt10m_y_2d:units = "m s-1" ;
		Mesh2_face_WindVelocityAt10m_y_2d:mesh = "Mesh2" ;
	float Mesh2_face_WindVelocityAt10m_x_2d(nMesh2_data_time, nMesh2_face) ;
		Mesh2_face_WindVelocityAt10m_x_2d:_FillValue = 1.e+31f ;
		Mesh2_face_WindVelocityAt10m_x_2d:grid_mapping = "Mesh2_crs" ;
		Mesh2_face_WindVelocityAt10m_x_2d:coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ;
		Mesh2_face_WindVelocityAt10m_x_2d:long_name = "wind_velocityAt10m (x-Komponente), Face (Polygon)" ;
		Mesh2_face_WindVelocityAt10m_x_2d:standard_name = "wind_x_velocityAt10m" ;
		Mesh2_face_WindVelocityAt10m_x_2d:cell_methods = "nMesh2_data_time: point nMesh2_layer_2d: mean area: point" ;
		Mesh2_face_WindVelocityAt10m_x_2d:name_id = 557 ;
		Mesh2_face_WindVelocityAt10m_x_2d:location = "face" ;
		Mesh2_face_WindVelocityAt10m_x_2d:units = "m s-1" ;
		Mesh2_face_WindVelocityAt10m_x_2d:mesh = "Mesh2" ;

// global attributes:
		:title = "mossco >>> uGrid conversion" ;
		:history = "Createded on Fri Jun 26 16:48:33 2015" ;
		:Conventions = "CF-1.6" ;
		:references = "http://www.baw.de/ und http://www.baw.de/methoden/index.php5/NetCDF" ;
}
