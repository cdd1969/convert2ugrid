float Mesh2_face_Stroemungsgeschwindigkeit_x_2d(nMesh2_data_time, nMesh2_layer_2d, nMesh2_face) ;
    Mesh2_face_Stroemungsgeschwindigkeit_x_2d:long_name = "Stroemungsgeschwindigkeit (x-Komponente), Face (Polygon)" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_x_2d:units = "m s-1" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_x_2d:name_id = 2 ; 
    Mesh2_face_Stroemungsgeschwindigkeit_x_2d:_FillValue = 1.e+31f ; 
    Mesh2_face_Stroemungsgeschwindigkeit_x_2d:cell_methods = "nMesh2_data_time: point nMesh2_layer_2d: mean area: point" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_x_2d:coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat Mesh2_face_z_face_2d" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_x_2d:grid_mapping = "Mesh2_crs" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_x_2d:standard_name = "sea_water_x_velocity" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_x_2d:mesh = "Mesh2" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_x_2d:location = "face" ; 
//    Mesh2_face_Stroemungsgeschwindigkeit_x_2d:davit_role = "visualization_variable" ;



float Mesh2_face_Stroemungsgeschwindigkeit_y_2d(nMesh2_data_time, nMesh2_layer_2d, nMesh2_face) ;
    Mesh2_face_Stroemungsgeschwindigkeit_y_2d:long_name = "Stroemungsgeschwindigkeit (y-Komponente), Face (Polygon)" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_y_2d:units = "m s-1" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_y_2d:name_id = 2 ; 
    Mesh2_face_Stroemungsgeschwindigkeit_y_2d:_FillValue = 1.e+31f ; 
    Mesh2_face_Stroemungsgeschwindigkeit_y_2d:cell_methods = "nMesh2_data_time: point nMesh2_layer_2d: mean area: point" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_y_2d:coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat Mesh2_face_z_face_2d" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_y_2d:grid_mapping = "Mesh2_crs" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_y_2d:standard_name = "sea_water_y_velocity" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_y_2d:mesh = "Mesh2" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_y_2d:location = "face" ; 
//    Mesh2_face_Stroemungsgeschwindigkeit_y_2d:davit_role = "visualization_variable" ;


float Mesh2_face_Stroemungsgeschwindigkeit_m_2d(nMesh2_data_time, nMesh2_layer_2d, nMesh2_face) ;
    Mesh2_face_Stroemungsgeschwindigkeit_m_2d:long_name = "Stroemungsgeschwindigkeit (Betrag), Face (Polygon)" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_m_2d:units = "m s-1" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_m_2d:name_id = 2 ; 
    Mesh2_face_Stroemungsgeschwindigkeit_m_2d:_FillValue = 1.e+31f ; 
    Mesh2_face_Stroemungsgeschwindigkeit_m_2d:cell_methods = "nMesh2_data_time: point nMesh2_layer_2d: mean area: point" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_m_2d:coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat Mesh2_face_z_face_2d" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_m_2d:grid_mapping = "Mesh2_crs" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_m_2d:standard_name = "magnitude_of_sea_water_velocity" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_m_2d:mesh = "Mesh2" ; 
    Mesh2_face_Stroemungsgeschwindigkeit_m_2d:location = "face" ; 
//    Mesh2_face_Stroemungsgeschwindigkeit_m_2d:davit_role = "visualization_variable" ;

   
float Mesh2_face_Temperatur_3d(nMesh2_data_time, nMesh2_layer_3d, nMesh2_face) ;
    Mesh2_face_Temperatur_3d:long_name = "Temperatur, Face (Polygon)" ;
    Mesh2_face_Temperatur_3d:units = "degC" ;
    Mesh2_face_Temperatur_3d:name_id = 6 ;
    Mesh2_face_Temperatur_3d:_FillValue = 1.e+31f ;
    Mesh2_face_Temperatur_3d:cell_measures = "area: Mesh2_face_wet_area" ;
    Mesh2_face_Temperatur_3d:cell_methods = "nMesh2_data_time: point nMesh2_layer_3d: mean area: point" ;
    Mesh2_face_Temperatur_3d:coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat Mesh2_face_z_face_3d" ;
    Mesh2_face_Temperatur_3d:grid_mapping = "Mesh2_crs" ;
    Mesh2_face_Temperatur_3d:standard_name = "temperature" ;
    Mesh2_face_Temperatur_3d:mesh = "Mesh2" ;
    Mesh2_face_Temperatur_3d:location = "face" ;
//    Mesh2_face_Temperatur_3d:davit_role = "visualization_variable" ;

double Mesh2_face_depth_2d(nMesh2_time, nMesh2_face) ;
    Mesh2_face_depth_2d:long_name = "Topographie" ;
    Mesh2_face_depth_2d:units = "m" ;
    Mesh2_face_depth_2d:name_id = 17 ;
    Mesh2_face_depth_2d:valid_range = -8848., 11034. ;
    Mesh2_face_depth_2d:_FillValue = 1.e+31 ;
    Mesh2_face_depth_2d:cell_measures = "area: Mesh2_face_area" ;
    Mesh2_face_depth_2d:cell_methods = "nMesh2_time: mean area: mean" ;
    Mesh2_face_depth_2d:coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ;
    Mesh2_face_depth_2d:grid_mapping = "Mesh2_crs" ;
    Mesh2_face_depth_2d:standard_name = "sea_floor_depth_below_geoid" ;
    Mesh2_face_depth_2d:mesh = "Mesh2" ;
    Mesh2_face_depth_2d:location = "face" ;
//    Mesh2_face_depth_2d:davit_role = "visualization_variable" ;

float Mesh2_face_Wasserstand_2d(nMesh2_data_time, nMesh2_face) ;
    Mesh2_face_Wasserstand_2d:long_name = "Wasserstand, Face (Polygon)" ; 
    Mesh2_face_Wasserstand_2d:units = "m" ; 
    Mesh2_face_Wasserstand_2d:name_id = 3 ; 
    Mesh2_face_Wasserstand_2d:_FillValue = 1.e+31f ; 
    Mesh2_face_Wasserstand_2d:cell_measures = "area: Mesh2_face_wet_area" ; 
    Mesh2_face_Wasserstand_2d:cell_methods = "nMesh2_data_time: point area: mean" ; 
    Mesh2_face_Wasserstand_2d:coordinates = "Mesh2_face_x Mesh2_face_y Mesh2_face_lon Mesh2_face_lat" ; 
    Mesh2_face_Wasserstand_2d:grid_mapping = "Mesh2_crs" ; 
    Mesh2_face_Wasserstand_2d:standard_name = "sea_surface_height" ; 
    Mesh2_face_Wasserstand_2d:mesh = "Mesh2" ; 
    Mesh2_face_Wasserstand_2d:location = "face" ; 

float Mesh2_face_Gesamtwassertiefe_2d(nMesh2_data_time, nMesh2_face) ;
    Mesh2_face_Gesamtwassertiefe_2d:long_name = "Gesamtwassertiefe [ face ]" ;
    Mesh2_face_Gesamtwassertiefe_2d:units = "m" ;
    Mesh2_face_Gesamtwassertiefe_2d:name_id = 16 ;
    Mesh2_face_Gesamtwassertiefe_2d:_FillValue = 1.e+31f ;
    Mesh2_face_Gesamtwassertiefe_2d:cell_methods = "nMesh2_data_time: point nMesh2_face: mean" ;
    Mesh2_face_Gesamtwassertiefe_2d:coordinates = "Mesh2_face_lon Mesh2_face_lat Mesh2_face_x Mesh2_face_y" ;
    Mesh2_face_Gesamtwassertiefe_2d:grid_mapping = "Mesh2_crs" ;
    Mesh2_face_Gesamtwassertiefe_2d:standard_name = "sea_floor_depth_below_sea_surface" ;
    Mesh2_face_Gesamtwassertiefe_2d:mesh = "Mesh2" ;
    Mesh2_face_Gesamtwassertiefe_2d:location = "face" ;
